module testClock;
    parameter WIDTH = 8;

    output [WIDTH-1 : 0] out;
    input clk, reset;

    reg [WIDTH-1 : 0] out;
    wire clk, reset;

    
endmodule